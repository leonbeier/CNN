library ieee;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;
    
library work;
    use work.bitwidths.all;
    use work.cnn_types.all;
    
entity multi_conv_comb is
    generic(
        PIXEL_SIZE: integer := 8;
        IMAGE_WIDTH: integer := 28
        
    );
    port(
    clk: in std_logic;
    reset_n: in std_logic;
    enable: in std_logic;
    in_data: in std_logic_vector(PIXEL_SIZE-1 downto 0);
    in_dv: in std_logic;
    in_fv: in std_logic;
    -- Reduce the I/O
    --out_data      : out final_pixel_array (9 downto 0);
    prediction    : out std_logic_vector (3 downto 0);
    out_fv        : out std_logic ;
    out_step_warning : out std_logic
    );
end entity;


architecture STRUCTURAL of multi_conv_comb is
constant  CONV1_KERNEL_VALUE_1 : 
            pixel_array := ("00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111","00000111");
constant  CONV1_KERNEL_VALUE_2 : 
        pixel_array := ("11100001","11100001","11100001","11100001","11100001","11100001","11100001","11100001","11100001");
        
--constant  CONV1_KERNEL_VALUE_1 : 
--            pixel_array := ("01001001","00011110","00000000","11110101","11111111","10110001","11000110","11100110","11000110");
--constant  CONV1_KERNEL_VALUE_2 : 
--        pixel_array := ("00011000","01011101","11001100","00110000","11100100","11111001","00100110","11010110","11101000");



constant CONV1_BIAS_VALUE_1 :
                        std_logic_vector := ("00000000");
 
constant CONV1_BIAS_VALUE_2 :
                        std_logic_vector := ("00000000");
--constant CONV1_BIAS_VALUE_3 :
--                        std_logic_vector := ("00000");
                        


constant MY_INT_MATRIX :
        int_matrix := ((233,230,169,160,169,205,208,168,151,170),(218,236,184,164,170,207,211,176,156,169),(206,167,195,210,143,218,218,165,150,164),(194,162,184,224,142,208,219,174,150,167),(167,129,201,203,158,136,231,140,88,160),(174,143,208,208,168,136,227,146,119,176),(176,166,219,197,143,170,221,117,146,137),(175,180,220,203,165,187,226,130,166,141),(179,177,216,201,172,183,219,106,169,94),(185,175,209,200,182,186,225,119,173,116),(189,188,210,201,166,179,211,105,171,55),(188,204,207,201,179,185,216,118,172,84),(180,202,202,199,184,186,206,108,177,66),(180,211,201,196,190,192,212,123,173,81),(183,200,206,201,183,196,207,116,183,95),(191,202,199,199,189,192,215,142,189,118),(182,179,201,199,169,199,210,129,176,169),(185,180,193,193,180,197,218,145,174,187),(179,171,189,197,174,205,217,156,168,133),(186,169,176,176,204,191,226,139,170,117),(175,157,195,171,185,200,229,149,182,148),(186,174,189,124,210,174,238,161,196,162),(167,130,218,126,152,181,232,177,171,167),(181,143,227,143,152,166,226,178,158,179),(177,157,233,180,144,196,204,191,146,183),(181,160,195,183,165,212,215,196,152,192),(200,229,187,215,163,181,192,200,211,169),(221,243,199,212,156,192,178,194,187,155),(157,229,189,213,200,166,213,191,147,137),(156,220,195,208,203,170,210,193,160,133),(182,200,199,207,203,189,190,190,188,120),(186,200,203,206,202,188,199,194,194,131),(197,196,205,205,199,192,192,191,196,152),(193,197,200,204,206,192,202,189,197,162),(198,202,205,205,195,195,191,180,201,186),(199,207,203,203,202,196,203,174,198,185),(200,203,207,206,195,197,192,185,204,194),(206,210,205,201,207,196,206,185,207,188),(202,199,207,206,192,197,194,184,204,193),(207,211,201,199,205,196,208,164,208,172),(205,201,207,206,191,203,201,188,207,192),(208,211,197,195,206,199,213,169,209,164),(204,195,204,202,189,205,203,169,206,188),(207,215,188,181,211,201,219,162,207,168),(202,195,199,199,189,207,207,144,204,183),(198,218,161,159,221,204,222,140,207,158),(199,199,196,192,192,207,210,152,202,163),(209,219,153,166,218,206,218,171,197,114),(197,195,179,179,200,214,224,101,194,62),(184,181,174,101,208,207,224,88,195,82),(180,144,173,55,193,223,218,133,197,107),(146,150,155,141,172,220,221,152,216,147),(149,189,197,219,178,192,185,225,104,121),(164,189,206,214,193,181,161,221,109,124),(188,195,201,211,203,174,194,210,191,126),(193,202,199,205,204,188,199,202,194,138),(193,196,202,206,203,191,185,207,197,180),(197,188,201,206,203,198,204,210,201,184),(191,189,203,207,203,197,185,208,200,196),(195,189,201,201,209,197,204,206,202,195),(199,192,203,207,202,200,185,206,203,201),(200,198,201,199,206,198,201,203,204,198),(202,196,206,208,198,203,190,204,207,206),(201,199,198,196,202,196,202,191,203,199),(202,192,201,204,188,197,187,198,203,204),(205,203,199,190,204,198,207,184,205,201),(204,194,203,204,186,201,189,198,204,205),(208,207,192,184,216,193,210,190,203,195),(204,191,200,201,191,202,185,199,205,204),(206,216,180,172,225,194,209,198,203,185),(204,193,198,201,195,206,189,199,207,202),(200,218,164,156,224,201,196,196,201,177),(202,197,195,195,197,209,201,195,205,196),(195,227,167,145,229,205,193,190,204,170),(199,197,183,179,200,211,214,182,203,172),(155,208,163,52,231,210,202,176,214,130),(161,166,138,102,202,230,228,115,201,132),(162,142,171,98,208,220,207,115,199,103),(218,181,203,206,195,104,146,222,196,147),(204,180,202,201,192,122,161,211,201,169),(181,206,198,211,200,164,159,216,203,186),(197,179,196,202,202,193,198,202,200,191),(194,195,202,205,194,186,180,212,199,196),(201,186,199,201,201,198,207,203,203,198),(198,198,199,204,197,192,182,208,199,197),(203,185,199,199,204,200,207,203,205,201),(197,188,203,205,195,194,182,208,203,202),(205,196,200,194,207,202,205,202,207,204),(199,180,205,206,194,199,183,208,205,206),(202,198,194,191,206,199,203,195,203,205),(203,190,206,204,188,199,185,209,203,209),(202,199,196,194,207,192,204,184,199,200),(208,194,205,204,184,202,182,208,202,207),(208,206,204,198,224,183,200,193,200,196),(210,180,200,202,192,202,185,206,203,207),(196,209,205,198,223,174,192,194,205,189),(208,169,194,196,195,204,196,203,205,202),(194,205,204,193,225,172,197,199,205,189),(209,178,191,193,201,209,209,203,211,200),(190,204,200,189,222,187,174,205,204,182),(206,184,179,182,197,214,202,194,211,188),(173,149,191,94,225,199,187,208,205,163),(187,149,107,49,209,243,186,173,217,159),(146,173,159,173,191,209,195,213,213,73),(224,194,195,212,178,100,147,224,151,172),(212,180,198,202,196,101,162,204,195,188),(191,181,206,209,183,192,164,211,193,193),(200,179,192,196,199,202,202,198,201,203),(207,197,212,209,193,188,190,209,195,199),(207,192,191,193,201,202,207,196,203,203),(204,208,204,204,203,190,188,211,202,204),(203,184,189,187,204,200,205,196,204,204),(197,202,194,204,204,194,178,209,206,207),(206,194,193,192,210,202,206,197,205,207),(193,186,195,208,198,201,182,210,209,205),(199,197,183,198,208,196,202,187,200,202),(187,201,193,207,188,208,187,209,212,195),(197,204,196,205,206,183,200,194,198,203),(183,205,194,203,185,209,196,205,204,198),(200,203,208,206,218,163,192,202,206,208),(196,175,193,201,197,209,203,202,202,206),(206,185,210,203,216,129,194,201,209,209),(203,171,190,192,199,203,208,200,209,206),(207,171,210,195,214,117,188,194,207,201),(211,175,188,176,201,203,216,200,209,203),(216,219,215,187,212,124,175,202,214,202),(215,195,187,176,197,208,219,194,212,187),(220,208,229,181,204,145,162,177,209,185),(181,182,157,56,186,242,194,163,223,154),(155,251,220,236,167,191,188,185,199,156),(201,206,163,180,173,197,140,237,207,177),(192,187,181,193,205,194,139,205,189,202),(208,209,211,208,188,170,169,220,189,194),(210,193,184,184,203,201,208,201,202,212),(208,200,212,209,207,177,190,209,184,195),(210,186,179,180,207,203,208,197,200,207),(201,206,200,210,209,188,187,211,197,198),(206,192,183,193,209,202,210,198,200,208),(197,193,201,214,205,201,183,196,208,203),(206,192,184,204,210,202,207,194,201,207),(177,188,203,211,204,209,181,182,212,207),(198,202,188,208,203,196,204,176,200,198),(158,186,200,206,205,211,199,176,210,209),(177,205,198,205,197,176,195,202,195,205),(151,195,192,202,199,211,211,184,208,207),(203,195,207,199,211,142,199,213,203,206),(169,178,182,204,200,212,211,192,206,210),(213,170,213,190,208,112,194,212,206,204),(191,168,184,201,202,206,211,194,201,205),(218,216,215,169,211,104,200,204,208,204),(203,179,189,192,210,200,215,197,202,201),(220,212,215,159,205,80,211,192,211,201),(217,195,200,165,207,186,224,197,204,191),(215,213,237,208,206,107,203,156,173,204),(204,175,219,122,184,207,199,159,214,134),(194,226,250,222,165,160,168,164,123,192),(174,231,194,205,197,162,133,233,160,151),(177,227,186,186,215,198,136,205,205,210),(213,205,221,220,210,177,153,209,146,173),(212,213,178,178,208,195,209,199,188,207),(202,180,227,215,204,181,186,202,190,184),(209,185,183,180,208,195,208,197,187,205),(199,201,218,208,198,188,182,196,202,200),(209,193,193,197,208,198,210,195,194,204),(184,194,210,206,198,195,179,190,206,207),(204,187,194,204,202,198,207,189,196,200),(165,187,209,205,210,206,188,187,205,211),(192,210,204,210,182,194,204,189,205,190),(165,164,208,201,210,214,214,183,203,208),(177,211,207,205,196,184,207,214,196,205),(169,191,201,202,197,211,215,176,201,199),(208,192,208,189,206,176,207,216,199,202),(172,175,188,204,200,206,212,196,200,191),(212,191,207,181,200,181,192,213,188,197),(182,155,192,206,210,203,211,211,199,191),(211,210,210,179,203,174,206,207,178,204),(191,160,195,198,210,199,206,210,194,184),(217,209,203,155,200,167,213,203,166,205),(207,194,206,187,206,194,210,202,190,173),(212,182,218,164,197,156,211,166,177,188),(217,208,231,150,204,174,212,191,187,126),(149,222,244,194,190,122,157,182,114,212),(159,233,216,232,190,178,132,216,185,137),(160,218,208,209,203,187,134,191,190,207),(205,191,213,217,192,211,151,200,175,166),(211,179,201,192,202,188,207,197,179,198),(186,183,216,215,194,215,172,199,209,185),(212,176,203,185,207,190,210,198,195,201),(179,188,209,202,187,199,174,200,207,203),(211,187,204,190,205,190,210,196,201,201),(182,194,206,199,202,195,181,200,203,216),(203,195,204,190,189,189,206,195,204,186),(187,171,208,197,209,205,196,200,197,216),(185,209,208,198,178,191,208,204,210,183),(189,147,209,201,209,210,213,192,193,206),(195,207,205,189,195,192,213,211,194,200),(199,185,204,206,198,211,215,187,205,191),(208,181,200,195,201,196,205,216,185,204),(189,181,196,207,201,206,208,198,207,177),(211,185,200,199,197,201,204,216,180,202),(184,175,201,206,208,201,205,205,202,180),(209,197,194,191,194,196,207,209,176,199),(181,187,210,199,207,198,199,203,200,181),(214,189,190,193,188,202,215,206,187,203),(200,205,213,189,205,192,197,190,197,173),(207,209,194,164,168,213,212,162,192,175),(207,208,231,168,201,175,214,164,181,89),(165,204,242,178,215,112,151,162,112,194),(160,187,212,224,201,186,152,226,135,144),(189,187,215,219,194,187,149,200,161,194),(182,122,216,222,213,213,147,196,199,141),(209,156,208,202,193,191,197,196,195,190),(175,191,213,223,185,218,154,188,201,198),(211,193,210,196,201,194,205,196,205,194),(181,198,208,215,175,215,178,195,202,202),(206,198,208,187,193,187,205,198,207,187),(194,185,199,212,190,212,186,195,196,215),(204,203,209,183,191,189,208,202,213,185),(204,162,198,210,201,209,199,197,181,215),(191,207,209,185,197,191,201,204,210,195),(209,160,206,214,204,205,208,194,185,201),(198,202,197,192,201,193,203,203,195,201),(205,188,206,212,186,206,210,177,208,175),(209,178,199,205,204,201,206,205,198,205),(198,201,208,207,190,204,210,192,211,159),(206,183,188,200,194,201,204,200,191,199),(188,206,212,201,195,195,204,198,205,179),(213,190,191,201,193,204,206,200,197,202),(179,214,216,193,204,199,200,190,200,193),(216,170,185,208,180,210,207,170,200,200),(188,209,221,186,204,200,195,180,200,194),(203,201,175,195,177,209,208,194,196,210),(198,222,233,129,190,197,203,181,183,141),(196,224,208,130,200,135,196,186,128,202),(199,206,204,212,171,197,125,224,162,106),(207,197,217,216,188,184,141,193,170,184),(159,215,208,221,175,212,146,183,185,191),(211,199,213,207,187,192,189,196,204,191),(175,218,205,226,162,223,147,190,193,191),(204,200,209,202,180,196,194,190,206,186),(185,205,198,216,176,216,179,197,187,208),(204,203,210,198,187,196,200,199,209,190),(202,202,197,213,180,215,192,197,188,205),(201,201,204,190,196,194,200,200,207,193),(207,197,197,213,172,210,200,192,196,204),(191,202,198,192,203,193,192,205,205,201),(211,181,202,213,154,209,208,178,203,193),(196,200,189,202,207,197,181,205,203,205),(210,194,207,207,165,206,208,165,206,168),(202,181,192,202,205,201,194,199,202,205),(204,214,215,205,184,207,209,164,210,165),(205,165,186,202,202,204,200,196,202,203),(194,213,219,196,196,199,206,169,203,192),(209,152,185,201,199,207,197,188,205,204),(182,213,222,187,208,198,202,168,199,204),(209,151,178,198,185,210,186,183,206,200),(178,206,224,182,210,203,195,145,204,212),(174,211,167,186,188,210,190,219,200,236),(183,229,231,110,176,199,186,181,159,202),(230,228,178,198,193,160,219,204,123,182),(169,210,204,228,143,181,156,158,163,184),(195,206,219,206,168,168,142,128,177,182),(150,233,189,220,149,211,102,224,158,178),(208,210,212,205,148,187,135,212,203,195),(179,213,193,225,190,221,141,215,170,205),(202,205,208,205,182,194,174,208,204,194),(191,203,196,218,196,216,161,208,191,214),(198,201,204,204,194,200,187,206,202,200),(198,180,197,215,173,212,188,200,203,207),(198,201,199,199,199,201,194,208,202,203),(204,172,198,212,149,211,199,181,207,203),(184,204,190,200,205,202,194,209,206,206),(209,179,201,209,136,210,205,177,209,201),(183,207,183,200,208,202,164,206,205,205),(206,195,198,205,165,206,205,188,206,192),(185,202,192,201,209,202,169,201,205,208),(200,207,208,197,190,203,204,190,204,190),(180,210,193,199,208,200,178,194,203,205),(178,215,219,188,208,199,199,176,201,198),(196,177,189,198,208,206,185,189,205,207),(163,220,226,160,216,182,184,185,201,219),(179,187,185,196,206,209,185,198,204,206),(193,179,228,141,222,200,172,125,205,224),(156,218,180,191,192,208,180,204,204,236),(195,230,222,96,206,199,150,173,149,216),(244,255,176,224,198,165,218,153,146,162),(165,156,121,223,161,232,178,238,154,120),(137,153,204,214,141,204,171,212,173,182),(146,173,143,231,202,223,149,226,101,203),(194,207,201,203,161,177,59,219,191,203),(149,180,158,228,195,222,101,209,157,214),(191,204,200,206,201,185,119,219,196,205),(183,172,172,223,165,222,134,197,198,196),(182,201,193,205,198,196,142,208,191,203),(208,165,188,223,139,221,193,183,213,194),(189,203,189,209,204,202,157,211,197,207),(213,168,194,218,151,220,191,170,213,188),(174,206,181,206,201,202,172,208,198,207),(215,177,197,212,166,213,197,184,210,187),(142,213,165,201,208,199,153,208,194,208),(212,190,204,207,179,210,192,184,210,189),(133,218,189,203,214,203,97,206,190,212),(204,206,216,193,201,200,193,190,208,206),(154,231,187,198,210,200,121,192,188,209),(148,208,223,174,211,180,178,193,201,220),(151,224,188,207,206,210,160,192,193,210),(135,209,222,144,215,155,179,192,192,223),(163,209,177,206,205,219,139,203,190,205),(184,183,211,162,215,190,177,152,196,228),(175,201,173,220,199,220,151,205,190,196),(166,211,228,184,203,177,126,156,158,203),(188,248,197,205,235,148,208,153,144,179),(171,181,168,165,169,188,195,206,172,216),(160,138,122,195,166,229,187,245,144,163),(140,178,138,189,218,228,183,179,116,226),(141,159,103,216,218,147,138,214,131,225),(134,153,128,232,204,229,167,196,132,211),(144,185,131,222,199,161,77,226,167,223),(159,153,159,241,146,225,150,199,189,197),(138,189,79,220,200,186,0,225,161,217),(175,182,169,242,159,230,184,190,207,169),(124,156,98,215,200,200,84,217,174,214),(178,173,169,241,173,241,194,189,204,172),(127,187,87,212,189,200,140,213,185,210),(147,177,201,234,183,233,168,204,173,192),(94,175,119,201,194,192,103,213,181,209),(136,188,194,197,195,233,110,205,195,204),(120,172,109,211,193,204,94,213,176,217),(128,150,211,194,196,204,140,210,211,209),(83,175,114,213,192,201,70,209,173,222),(127,140,200,169,184,196,140,215,202,218),(115,182,145,210,171,211,104,208,159,228),(134,163,195,144,181,197,128,224,183,218),(142,165,140,130,189,234,154,221,179,192),(144,172,169,161,204,209,154,210,168,210),(171,193,180,169,220,222,175,212,156,189),(179,191,200,162,167,224,178,172,140,213),(194,203,192,183,182,186,198,217,183,188));
constant MY_INT_MATRIX_BIAS :
        int_array :=(63,255,92,73,93,140,74,139,0,82);



-- COMPONENTS
component firstLayer is
    generic(
    PIXEL_SIZE    :   integer ;
    IMAGE_WIDTH   :   integer ;
    KERNEL_SIZE   :   integer ;
    KERNEL_VALUE_1  :   pixel_array;
    KERNEL_VALUE_2  :   pixel_array;
--    KERNEL_VALUE_3  :   pixel_array;
    NB_IN_FLOWS   :   integer ;
    NB_OUT_FLOWS  :   integer ;
    BIAS_VALUE_1    :   std_logic_vector;
    BIAS_VALUE_2    :   std_logic_vector
--    BIAS_VALUE_3    :   std_logic_vector
);

port(
    clk           :   in  std_logic;
    reset_n       :   in  std_logic;
    enable        :   in  std_logic;
    in_data       :   in  std_logic_vector (PIXEL_SIZE-1 downto 0);
    in_dv         :   in  std_logic;
    in_fv         :   in  std_logic;

    out_data      :   out no_a_pixel_array (NB_OUT_FLOWS - 1 downto 0);
    out_dv        :   out std_logic_vector (NB_OUT_FLOWS - 1 downto 0);
    out_fv        :   out std_logic_vector (NB_OUT_FLOWS - 1 downto 0)
);
  end component;


  component poolLayer is
     generic(
     PIXEL_SIZE    :   integer;
     IMAGE_WIDTH   :   integer;
     KERNEL_SIZE   :   integer;
     NB_OUT_FLOWS  :   integer
 );

     port(
       clk           : in  std_logic;
       reset_n       : in  std_logic;
       enable        : in  std_logic;
       in_data       : in  no_a_pixel_array (0 to NB_OUT_FLOWS - 1);
       in_dv         : in  std_logic_vector (0 to NB_OUT_FLOWS - 1);
       in_fv         : in  std_logic_vector (0 to NB_OUT_FLOWS - 1);
       out_data      : out no_a_pixel_array (0 to NB_OUT_FLOWS - 1);
       out_dv        : out std_logic_vector (0 to NB_OUT_FLOWS - 1);
       out_fv        : out std_logic_vector (0 to NB_OUT_FLOWS - 1)
   );
  end component;
  component dsp_layer is
   generic(
       MY_MATRIX     :   int_matrix;
       MY_MATRIX_BIAS :  int_array;
       IMAGE_WIDTH   :   integer ;
       NB_IN_FLOWS   :   integer 
   );
 
       port(
         clk           : in  std_logic;
         reset_n       : in  std_logic;
         enable        : in  std_logic;
         in_data       : in  no_a_pixel_array (0 to NB_IN_FLOWS - 1);
         in_dv         : in  std_logic_vector (0 to NB_IN_FLOWS - 1);
         in_fv         : in  std_logic_vector (0 to NB_IN_FLOWS - 1);
         out_data      : out final_pixel_array (9 downto 0);
         prediction    : out std_logic_vector (3 downto 0);
         out_fv        : out std_logic ;
         out_step_warning : out std_logic
     );
end component;

   -- SIGNALS
 
 
   signal conv1_data : no_a_pixel_array (0 to 1);
   signal conv1_dv : std_logic_vector(0 to 1);
   signal conv1_fv : std_logic_vector(0 to 1);
   signal dsp_data : no_a_pixel_array (0 to 1);
   signal dsp_fv   : std_logic_vector (0 to 1);
   signal dsp_dv   : std_logic_vector (0 to 1);


 
   -- STRUCTURAL DESCRIPTION
  -- Deleted:
          --KERNEL_VALUE_3 => CONV1_KERNEL_VALUE_3,
          --BIAS_VALUE_3 => CONV1_BIAS_VALUE_3
 begin
   conv1: firstLayer
     generic map(
       PIXEL_SIZE => PIXEL_SIZE,
       IMAGE_WIDTH => 28,
       KERNEL_SIZE => 3,
       NB_IN_FLOWS => 1,
       NB_OUT_FLOWS => 2,
       KERNEL_VALUE_1 => CONV1_KERNEL_VALUE_1,
       KERNEL_VALUE_2 => CONV1_KERNEL_VALUE_2,
       BIAS_VALUE_1 => CONV1_BIAS_VALUE_1,
       BIAS_VALUE_2 => CONV1_BIAS_VALUE_2

     )
     port map(
       clk => clk,
       reset_n => reset_n,
       enable => enable,
       in_data => in_data,
       in_dv => in_dv,
       in_fv => in_fv,
       out_data => conv1_data,
       out_dv => conv1_dv,
       out_fv => conv1_fv
     );
 
   pool1: poolLayer
     generic map(
       PIXEL_SIZE => PIXEL_SIZE,
       IMAGE_WIDTH => 26,
       KERNEL_SIZE => 2,
       NB_OUT_FLOWS => 2
     )
     port map(
       clk => clk,
       reset_n => reset_n,
       enable => enable,
       in_data => conv1_data,
       in_dv => conv1_dv,
       in_fv => conv1_fv,
       out_data => dsp_data,
       out_dv => dsp_dv,
       out_fv => dsp_fv
     );
     
     dsp_1: dsp_layer
     generic map(
        MY_MATRIX => MY_INT_MATRIX,
        MY_MATRIX_BIAS => MY_INT_MATRIX_BIAS,
        IMAGE_WIDTH => 13,
        NB_IN_FLOWS => 2
     )
     port map(
              clk  => clk,
              reset_n => reset_n,
              enable  => enable,
              in_data => dsp_data,
              in_dv   => dsp_dv,
              in_fv   => dsp_fv,
              out_data => open,
              prediction => prediction,
              out_fv  => out_fv,
              out_step_warning => out_step_warning 
       );

end architecture;
