library ieee;
    use    ieee.std_logic_1164.all;
    use    ieee.numeric_std.all;
library work;
    use work.bitwidths.all;

package    cnn_types is

    -- Types
        type     int_matrix is array (0 to 337,0 to 9) of integer;
        type     int_array is array (0 to 9) of integer;
        type     no_a_pixel_matrix is array (0 to 337,0 to 9) of std_logic_vector (SUM_WIDTH - 1 downto 0);
        type     no_a_pixel_array is array (natural range <>) of std_logic_vector (SUM_WIDTH - 1 downto 0);
        --type     final_pixel_array is array (natural range <>) of signed (2*SUM_WIDTH - 1 downto 0); 
        --CPU compatibility test
        type     final_pixel_array is array (natural range <>) of unsigned (63 downto 0);
        ---
        type     pixel_array    is array ( natural range <> ) of std_logic_vector (PIXEL_CONST-1 downto 0);
        type     sum_array      is array ( natural range <> ) of std_logic_vector (SUM_WIDTH-1 downto 0);
        type     pixel_matrix   is array ( natural range <> ,  natural range <>) of std_logic_vector (PIXEL_CONST-1 downto 0);
        
    ------------------------------------------------------------------------------

    -- Constants  : cf sumElement.vhd , TanH function ...
    constant SCALE_FACTOR      :   integer := 2 **(PIXEL_CONST-1) - 1;
    constant A1                :   integer := PIXEL_CONST - 1;
    constant A2                :   integer := PIXEL_CONST;
    constant T1                :   integer := SCALE_FACTOR * SCALE_FACTOR / 2;
    constant T2                :   integer := SCALE_FACTOR * SCALE_FACTOR * 5/4;
    constant V1                :   integer := SCALE_FACTOR / 4;
    constant V2                :   integer := SCALE_FACTOR - 10;

    ------------------------------------------------------------------------------

    -- Functions:
    -- extractRow : Extracts a row of pixel_array data from a pixel_matrix.
--    function extractRow( target_row :  integer;
--                            nb_col     :  integer;
--                            in_matrix  :  pixel_matrix )
--                            return        pixel_array;
--    ------------------------------------------------------------------------------
end cnn_types;


package body cnn_types is
--    function extractRow( target_row :  integer;
--                            nb_col     :  integer;
--                            in_matrix  :  pixel_matrix )
--                            return        pixel_array is
--    variable out_vec : pixel_array  (0 to nb_col - 1);
--    begin
--        for index_col in 0 to (nb_col - 1) loop
--            out_vec(index_col) := in_matrix(target_row,index_col);
--        end loop;
--        return out_vec;
--    end extractRow;

end cnn_types;